module tb_risc;

  reg clk;
  
  reg reset;
  
  risc dut(clk, reset);
  
  initial begin
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
     clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
     clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
        clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
    clk = 0;
    #5;
    clk = 1;
    #5;
  end
  
  initial begin
    reset = 1;
    repeat(5) @(posedge clk);
    reset = 0;
    #400;
    $finish;
  end
  
endmodule